library ieee;
use ieee.std_logic_1164.all; -- 1
-- 2
use ieee.numeric_std.all; /* 3 */

entity test2800 is
end test2800;

/* 4
5 
6*/