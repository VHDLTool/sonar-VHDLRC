package b is
  use c.all;
end;