-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés

library
print("Hello world")
print("Bonjour tout le monde")

-- Commentaire en français
-- Commentaire en français
-- Commentaire en français