 -- buffer
 -- Creation date
 -- License : Linty
 
 library IEEE;
 use IEEE.STD_LOGIC_1164.ALL;
 
 ENTITY test4200 IS
 end test4200;