an other line