library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY test2600 IS
 Port ( a : in std_logic;
 b : in std_logic;
 c : in std_logic;
 s : out std_logic);
end test2600;