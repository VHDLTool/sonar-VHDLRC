type test_type is array (0 to 7) of std_logic_vector(7 downto 0);
type test_type_issue is array (7 downto 0) of std_logic_vector(0 to 7);