-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés

library
hello

-- Commentaire en français
-- Commentaire en français
-- Commentaire en français
-- Commentaire en français

code

-- english comment

code

/*commentaire en
francais commentaire en
francais commentaire en
francais commentaire en
francais*/

code

-- commentaire commentaire commentaire commentaire commentaire commentaire commentaire commentaire commentaire commentaire

code

-- commentaire trop court

code

-- Demain tomorrow Demain tomorrow Demain tomorrow Demain tomorrow Demain tomorrow

code

-- Commentaire en français
-- Commentaire en français
-- Commentaire en français
-- Commentaire en français