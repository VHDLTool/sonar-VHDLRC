package d is
  use e.all;
end;