-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés

library
hello

-- Commentaire en français
-- Commentaire en français

code

/*commentaire en
francais*/

code

-- commentaire

code

-- commentaire non fiable ahghujhukjjklmkmlkklm

code

-- Commentaire en français
-- Commentaire en français