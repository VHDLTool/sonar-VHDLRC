-- entity hello_world is
-- end;
