package c is
  use d.all;
end;