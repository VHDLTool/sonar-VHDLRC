-- English header. All rights reserved
-- En-tête français. Tous drois réservés

print("Hello world")
print("Bonjour tout le monde")