-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés
-- En-tête français. Tous droits réservés

library
hello

-- English comment
-- English comment
-- English comment
-- English comment
-- English comment

code

-- Commentaire en français
-- Commentaire en français
-- Commentaire en français
-- Commentaire en français