library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY test2000 IS
    Port ( a : in std_logic; -- Indented with 4 spaces
    b : in std_logic; -- Indented with 4 spaces
	c : in std_logic; -- Indented with tab
    s : out std_logic); -- Indented with 4 spaces
end test2000;