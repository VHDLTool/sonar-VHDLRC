-------------------------------------------------------------------------------------------------
-- Author: Mickael Carl
-- Date: 2015-04-02
-------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;