package a is
  use b.all;
end;